module tb_top();
endmodule

module tb_top2();
endmodule
